---------------------------------------------------------------------------------------------------
-- Copyright (c) 2024 by XTools, Switzerland
---------------------------------------------------------------------------------------------------

---------------------------------------------------------------------------------------------------
-- Libraries
---------------------------------------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

library work;

---------------------------------------------------------------------------------------------------
-- Packet Header
---------------------------------------------------------------------------------------------------
package IpPackager_2020_1_pkg is

    -----------------------------------------------------------------------------------------------
    -- Constants
    -----------------------------------------------------------------------------------------------
    -- constant TestSlv_Width_c : integer := 2;
    constant TestSlv_Width_c : integer := integer(ceil(log2(real(3))));
    -- constant TestSlv_Width_c : integer := 2;

end package IpPackager_2020_1_pkg;


---------------------------------------------------------------------------------------------------
-- Packet Body
---------------------------------------------------------------------------------------------------
package body IpPackager_2020_1_pkg is

end package body IpPackager_2020_1_pkg;

---------------------------------------------------------------------------------------------------
-- EOF
---------------------------------------------------------------------------------------------------
